----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Kyara McWilliam
-- 
-- Create Date: 27.09.2024 10:47:43
-- Design Name: 
-- Module Name: Mux16_32bit_23375183 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Mux16_32bit_23375183 is
    Port (
        IN00, IN01, IN02, IN03, IN04, IN05, IN06, IN07, 
        IN08, IN09, IN10, IN11, IN12, IN13, IN14, IN15 : in STD_LOGIC_VECTOR (31 downto 0);
        S : in STD_LOGIC_VECTOR (3 downto 0); -- 4-bit selection signal
        Y : out STD_LOGIC_VECTOR (31 downto 0)
    );
end Mux16_32bit_23375183;

architecture Behavioral of Mux16_32bit_23375183 is

    -- 1-bit 16-input multiplexer component
    COMPONENT Mux16_1bit_23375183
        Port (
            I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15 : in STD_LOGIC;
            S : in STD_LOGIC_VECTOR (3 downto 0);
            Y : out STD_LOGIC
        );
    END COMPONENT;

begin

    -- For each bit of the output, instantiate a 1-bit 16-input multiplexer
    bit0: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(0), I1 => IN01(0), I2 => IN02(0), I3 => IN03(0),
        I4 => IN04(0), I5 => IN05(0), I6 => IN06(0), I7 => IN07(0),
        I8 => IN08(0), I9 => IN09(0), I10 => IN10(0), I11 => IN11(0),
        I12 => IN12(0), I13 => IN13(0), I14 => IN14(0), I15 => IN15(0),
        S => S,
        Y => Y(0)
    );

    bit1: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(1), I1 => IN01(1), I2 => IN02(1), I3 => IN03(1),
        I4 => IN04(1), I5 => IN05(1), I6 => IN06(1), I7 => IN07(1),
        I8 => IN08(1), I9 => IN09(1), I10 => IN10(1), I11 => IN11(1),
        I12 => IN12(1), I13 => IN13(1), I14 => IN14(1), I15 => IN15(1),
        S => S,
        Y => Y(1)
    );

    bit2: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(2), I1 => IN01(2), I2 => IN02(2), I3 => IN03(2),
        I4 => IN04(2), I5 => IN05(2), I6 => IN06(2), I7 => IN07(2),
        I8 => IN08(2), I9 => IN09(2), I10 => IN10(2), I11 => IN11(2),
        I12 => IN12(2), I13 => IN13(2), I14 => IN14(2), I15 => IN15(2),
        S => S,
        Y => Y(2)
    );

    bit3: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(3), I1 => IN01(3), I2 => IN02(3), I3 => IN03(3),
        I4 => IN04(3), I5 => IN05(3), I6 => IN06(3), I7 => IN07(3),
        I8 => IN08(3), I9 => IN09(3), I10 => IN10(3), I11 => IN11(3),
        I12 => IN12(3), I13 => IN13(3), I14 => IN14(3), I15 => IN15(3),
        S => S,
        Y => Y(3)
    );

    bit4: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(4), I1 => IN01(4), I2 => IN02(4), I3 => IN03(4),
        I4 => IN04(4), I5 => IN05(4), I6 => IN06(4), I7 => IN07(4),
        I8 => IN08(4), I9 => IN09(4), I10 => IN10(4), I11 => IN11(4),
        I12 => IN12(4), I13 => IN13(4), I14 => IN14(4), I15 => IN15(4),
        S => S,
        Y => Y(4)
    );

    bit5: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(5), I1 => IN01(5), I2 => IN02(5), I3 => IN03(5),
        I4 => IN04(5), I5 => IN05(5), I6 => IN06(5), I7 => IN07(5),
        I8 => IN08(5), I9 => IN09(5), I10 => IN10(5), I11 => IN11(5),
        I12 => IN12(5), I13 => IN13(5), I14 => IN14(5), I15 => IN15(5),
        S => S,
        Y => Y(5)
    );

    bit6: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(6), I1 => IN01(6), I2 => IN02(6), I3 => IN03(6),
        I4 => IN04(6), I5 => IN05(6), I6 => IN06(6), I7 => IN07(6),
        I8 => IN08(6), I9 => IN09(6), I10 => IN10(6), I11 => IN11(6),
        I12 => IN12(6), I13 => IN13(6), I14 => IN14(6), I15 => IN15(6),
        S => S,
        Y => Y(6)
    );

    bit7: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(7), I1 => IN01(7), I2 => IN02(7), I3 => IN03(7),
        I4 => IN04(7), I5 => IN05(7), I6 => IN06(7), I7 => IN07(7),
        I8 => IN08(7), I9 => IN09(7), I10 => IN10(7), I11 => IN11(7),
        I12 => IN12(7), I13 => IN13(7), I14 => IN14(7), I15 => IN15(7),
        S => S,
        Y => Y(7)
    );

    bit8: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(8), I1 => IN01(8), I2 => IN02(8), I3 => IN03(8),
        I4 => IN04(8), I5 => IN05(8), I6 => IN06(8), I7 => IN07(8),
        I8 => IN08(8), I9 => IN09(8), I10 => IN10(8), I11 => IN11(8),
        I12 => IN12(8), I13 => IN13(8), I14 => IN14(8), I15 => IN15(8),
        S => S,
        Y => Y(8)
    );

    bit9: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(9), I1 => IN01(9), I2 => IN02(9), I3 => IN03(9),
        I4 => IN04(9), I5 => IN05(9), I6 => IN06(9), I7 => IN07(9),
        I8 => IN08(9), I9 => IN09(9), I10 => IN10(9), I11 => IN11(9),
        I12 => IN12(9), I13 => IN13(9), I14 => IN14(9), I15 => IN15(9),
        S => S,
        Y => Y(9)
    );

    bit10: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(10), I1 => IN01(10), I2 => IN02(10), I3 => IN03(10),
        I4 => IN04(10), I5 => IN05(10), I6 => IN06(10), I7 => IN07(10),
        I8 => IN08(10), I9 => IN09(10), I10 => IN10(10), I11 => IN11(10),
        I12 => IN12(10), I13 => IN13(10), I14 => IN14(10), I15 => IN15(10),
        S => S,
        Y => Y(10)
    );

    bit11: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(11), I1 => IN01(11), I2 => IN02(11), I3 => IN03(11),
        I4 => IN04(11), I5 => IN05(11), I6 => IN06(11), I7 => IN07(11),
        I8 => IN08(11), I9 => IN09(11), I10 => IN10(11), I11 => IN11(11),
        I12 => IN12(11), I13 => IN13(11), I14 => IN14(11), I15 => IN15(11),
        S => S,
        Y => Y(11)
    );

    bit12: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(12), I1 => IN01(12), I2 => IN02(12), I3 => IN03(12),
        I4 => IN04(12), I5 => IN05(12), I6 => IN06(12), I7 => IN07(12),
        I8 => IN08(12), I9 => IN09(12), I10 => IN10(12), I11 => IN11(12),
        I12 => IN12(12), I13 => IN13(12), I14 => IN14(12), I15 => IN15(12),
        S => S,
        Y => Y(12)
    );

    bit13: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(13), I1 => IN01(13), I2 => IN02(13), I3 => IN03(13),
        I4 => IN04(13), I5 => IN05(13), I6 => IN06(13), I7 => IN07(13),
        I8 => IN08(13), I9 => IN09(13), I10 => IN10(13), I11 => IN11(13),
        I12 => IN12(13), I13 => IN13(13), I14 => IN14(13), I15 => IN15(13),
        S => S,
        Y => Y(13)
    );

    bit14: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(14), I1 => IN01(14), I2 => IN02(14), I3 => IN03(14),
        I4 => IN04(14), I5 => IN05(14), I6 => IN06(14), I7 => IN07(14),
        I8 => IN08(14), I9 => IN09(14), I10 => IN10(14), I11 => IN11(14),
        I12 => IN12(14), I13 => IN13(14), I14 => IN14(14), I15 => IN15(14),
        S => S,
        Y => Y(14)
    );

    bit15: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(15), I1 => IN01(15), I2 => IN02(15), I3 => IN03(15),
        I4 => IN04(15), I5 => IN05(15), I6 => IN06(15), I7 => IN07(15),
        I8 => IN08(15), I9 => IN09(15), I10 => IN10(15), I11 => IN11(15),
        I12 => IN12(15), I13 => IN13(15), I14 => IN14(15), I15 => IN15(15),
        S => S,
        Y => Y(15)
    );

    bit16: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(16), I1 => IN01(16), I2 => IN02(16), I3 => IN03(16),
        I4 => IN04(16), I5 => IN05(16), I6 => IN06(16), I7 => IN07(16),
        I8 => IN08(16), I9 => IN09(16), I10 => IN10(16), I11 => IN11(16),
        I12 => IN12(16), I13 => IN13(16), I14 => IN14(16), I15 => IN15(16),
        S => S,
        Y => Y(16)
    );

    bit17: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(17), I1 => IN01(17), I2 => IN02(17), I3 => IN03(17),
        I4 => IN04(17), I5 => IN05(17), I6 => IN06(17), I7 => IN07(17),
        I8 => IN08(17), I9 => IN09(17), I10 => IN10(17), I11 => IN11(17),
        I12 => IN12(17), I13 => IN13(17), I14 => IN14(17), I15 => IN15(17),
        S => S,
        Y => Y(17)
    );

    bit18: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(18), I1 => IN01(18), I2 => IN02(18), I3 => IN03(18),
        I4 => IN04(18), I5 => IN05(18), I6 => IN06(18), I7 => IN07(18),
        I8 => IN08(18), I9 => IN09(18), I10 => IN10(18), I11 => IN11(18),
        I12 => IN12(18), I13 => IN13(18), I14 => IN14(18), I15 => IN15(18),
        S => S,
        Y => Y(18)
    );

    bit19: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(19), I1 => IN01(19), I2 => IN02(19), I3 => IN03(19),
        I4 => IN04(19), I5 => IN05(19), I6 => IN06(19), I7 => IN07(19),
        I8 => IN08(19), I9 => IN09(19), I10 => IN10(19), I11 => IN11(19),
        I12 => IN12(19), I13 => IN13(19), I14 => IN14(19), I15 => IN15(19),
        S => S,
        Y => Y(19)
    );

    bit20: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(20), I1 => IN01(20), I2 => IN02(20), I3 => IN03(20),
        I4 => IN04(20), I5 => IN05(20), I6 => IN06(20), I7 => IN07(20),
        I8 => IN08(20), I9 => IN09(20), I10 => IN10(20), I11 => IN11(20),
        I12 => IN12(20), I13 => IN13(20), I14 => IN14(20), I15 => IN15(20),
        S => S,
        Y => Y(20)
    );

    bit21: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(21), I1 => IN01(21), I2 => IN02(21), I3 => IN03(21),
        I4 => IN04(21), I5 => IN05(21), I6 => IN06(21), I7 => IN07(21),
        I8 => IN08(21), I9 => IN09(21), I10 => IN10(21), I11 => IN11(21),
        I12 => IN12(21), I13 => IN13(21), I14 => IN14(21), I15 => IN15(21),
        S => S,
        Y => Y(21)
    );

    bit22: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(22), I1 => IN01(22), I2 => IN02(22), I3 => IN03(22),
        I4 => IN04(22), I5 => IN05(22), I6 => IN06(22), I7 => IN07(22),
        I8 => IN08(22), I9 => IN09(22), I10 => IN10(22), I11 => IN11(22),
        I12 => IN12(22), I13 => IN13(22), I14 => IN14(22), I15 => IN15(22),
        S => S,
        Y => Y(22)
    );

    bit23: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(23), I1 => IN01(23), I2 => IN02(23), I3 => IN03(23),
        I4 => IN04(23), I5 => IN05(23), I6 => IN06(23), I7 => IN07(23),
        I8 => IN08(23), I9 => IN09(23), I10 => IN10(23), I11 => IN11(23),
        I12 => IN12(23), I13 => IN13(23), I14 => IN14(23), I15 => IN15(23),
        S => S,
        Y => Y(23)
    );

    bit24: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(24), I1 => IN01(24), I2 => IN02(24), I3 => IN03(24),
        I4 => IN04(24), I5 => IN05(24), I6 => IN06(24), I7 => IN07(24),
        I8 => IN08(24), I9 => IN09(24), I10 => IN10(24), I11 => IN11(24),
        I12 => IN12(24), I13 => IN13(24), I14 => IN14(24), I15 => IN15(24),
        S => S,
        Y => Y(24)
    );

    bit25: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(25), I1 => IN01(25), I2 => IN02(25), I3 => IN03(25),
        I4 => IN04(25), I5 => IN05(25), I6 => IN06(25), I7 => IN07(25),
        I8 => IN08(25), I9 => IN09(25), I10 => IN10(25), I11 => IN11(25),
        I12 => IN12(25), I13 => IN13(25), I14 => IN14(25), I15 => IN15(25),
        S => S,
        Y => Y(25)
    );

    bit26: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(26), I1 => IN01(26), I2 => IN02(26), I3 => IN03(26),
        I4 => IN04(26), I5 => IN05(26), I6 => IN06(26), I7 => IN07(26),
        I8 => IN08(26), I9 => IN09(26), I10 => IN10(26), I11 => IN11(26),
        I12 => IN12(26), I13 => IN13(26), I14 => IN14(26), I15 => IN15(26),
        S => S,
        Y => Y(26)
    );

    bit27: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(27), I1 => IN01(27), I2 => IN02(27), I3 => IN03(27),
        I4 => IN04(27), I5 => IN05(27), I6 => IN06(27), I7 => IN07(27),
        I8 => IN08(27), I9 => IN09(27), I10 => IN10(27), I11 => IN11(27),
        I12 => IN12(27), I13 => IN13(27), I14 => IN14(27), I15 => IN15(27),
        S => S,
        Y => Y(27)
    );

    bit28: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(28), I1 => IN01(28), I2 => IN02(28), I3 => IN03(28),
        I4 => IN04(28), I5 => IN05(28), I6 => IN06(28), I7 => IN07(28),
        I8 => IN08(28), I9 => IN09(28), I10 => IN10(28), I11 => IN11(28),
        I12 => IN12(28), I13 => IN13(28), I14 => IN14(28), I15 => IN15(28),
        S => S,
        Y => Y(28)
    );

    bit29: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(29), I1 => IN01(29), I2 => IN02(29), I3 => IN03(29),
        I4 => IN04(29), I5 => IN05(29), I6 => IN06(29), I7 => IN07(29),
        I8 => IN08(29), I9 => IN09(29), I10 => IN10(29), I11 => IN11(29),
        I12 => IN12(29), I13 => IN13(29), I14 => IN14(29), I15 => IN15(29),
        S => S,
        Y => Y(29)
    );

    bit30: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(30), I1 => IN01(30), I2 => IN02(30), I3 => IN03(30),
        I4 => IN04(30), I5 => IN05(30), I6 => IN06(30), I7 => IN07(30),
        I8 => IN08(30), I9 => IN09(30), I10 => IN10(30), I11 => IN11(30),
        I12 => IN12(30), I13 => IN13(30), I14 => IN14(30), I15 => IN15(30),
        S => S,
        Y => Y(30)
    );

    bit31: Mux16_1bit_23375183 PORT MAP (
        I0 => IN00(31), I1 => IN01(31), I2 => IN02(31), I3 => IN03(31),
        I4 => IN04(31), I5 => IN05(31), I6 => IN06(31), I7 => IN07(31),
        I8 => IN08(31), I9 => IN09(31), I10 => IN10(31), I11 => IN11(31),
        I12 => IN12(31), I13 => IN13(31), I14 => IN14(31), I15 => IN15(31),
        S => S,
        Y => Y(31)
    );

end Behavioral;
